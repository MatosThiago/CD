library verilog;
use verilog.vl_types.all;
entity Coder is
    port(
        B0              : out    vl_logic;
        D1              : in     vl_logic;
        D5              : in     vl_logic;
        D9              : in     vl_logic;
        D7              : in     vl_logic;
        D3              : in     vl_logic;
        B1              : out    vl_logic;
        D2              : in     vl_logic;
        D6              : in     vl_logic;
        B2              : out    vl_logic;
        D4              : in     vl_logic;
        B3              : out    vl_logic;
        D8              : in     vl_logic;
        D0              : in     vl_logic
    );
end Coder;
