library verilog;
use verilog.vl_types.all;
entity Full_Adder_4_bits_vlg_vec_tst is
end Full_Adder_4_bits_vlg_vec_tst;
