library verilog;
use verilog.vl_types.all;
entity Subtractor_4_bits_vlg_vec_tst is
end Subtractor_4_bits_vlg_vec_tst;
