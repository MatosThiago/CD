library verilog;
use verilog.vl_types.all;
entity Subtractor_vlg_vec_tst is
end Subtractor_vlg_vec_tst;
