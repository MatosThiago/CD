library verilog;
use verilog.vl_types.all;
entity mux2_vlg_check_tst is
    port(
        F               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux2_vlg_check_tst;
