library verilog;
use verilog.vl_types.all;
entity Coder_vlg_vec_tst is
end Coder_vlg_vec_tst;
