library verilog;
use verilog.vl_types.all;
entity \4Bit_Multiplier\ is
    port(
        P0              : out    vl_logic;
        B0              : in     vl_logic;
        A0              : in     vl_logic;
        P1              : out    vl_logic;
        B1              : in     vl_logic;
        A1              : in     vl_logic;
        P2              : out    vl_logic;
        A2              : in     vl_logic;
        B2              : in     vl_logic;
        P3              : out    vl_logic;
        A3              : in     vl_logic;
        B3              : in     vl_logic;
        P4              : out    vl_logic;
        P5              : out    vl_logic;
        P6              : out    vl_logic;
        P7              : out    vl_logic
    );
end \4Bit_Multiplier\;
