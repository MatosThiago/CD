library verilog;
use verilog.vl_types.all;
entity Coder_vlg_check_tst is
    port(
        B0              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        B3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Coder_vlg_check_tst;
